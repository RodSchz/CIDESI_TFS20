* Netlist CIDESI_TFS10

.SUBCKT Resistor01
R$1 \$4 \$3 2.1528852459 RES1
R$2 \$6 \$5 3.83350819672 RES1
R$3 \$2 \$1 0.806596721311 RES1
.ENDS Resistor01
